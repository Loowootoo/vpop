/*
   中國古代數學家張丘建在他的《算經》
   提出了一個著名的「百錢買百雞問題」，
   雞翁一，值錢五，雞母一，值錢三，雞雛三，值錢一，
   百錢買百雞，問翁、母、雛各幾何？

   x = 翁
   y = 母
   z = 雛

   5x+3y+z/3 =100(百錢)
   x+y+z = 100(百雞)
   0 <= x <= 100/5 ==> range = 20
   0 <= y <= 100/3 ==> range = 33
   0 <= z <= 100   ==> range = 100
*/
module main

fn main() {
	mut x := 0
	mut y := 0
	mut z := 0
	mut sum := 0
	println("百錢買百雞問題")
	for x = 0; x <= 20; x++ {
		for y = 0; y <= 33; y++ {
			for z = 0; z <= 100; z++ {
				sum = 5 * x + 3 * y + z / 3
				if sum == 100 && z % 3 == 0 && x + y + z == 100 {
					println('翁:$x 母:$y 雛:$z')
				}
			}
		}
	}
}
